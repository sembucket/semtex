0.2  0.2  1.0  1.0
0.95 0.2  0.0  1.0
1.0  1.0  0.0  1.0
0.0  0.9  0.3  1.0
1.0  1.0  0.0  1.0
1.0  1.0  1.0  1.0
0.0  0.9  0.9  1.0
0.5  0.7  1.0  1.0
