# Example of a "script" for setting up an sview scene.
# Usage: sview -s tg.sv tg.mesh tg.fld

t 0 0.5 0
p -25 35 0
z 1.2
f u
m 0.4
a
f p
m -0.4
n
a
f w
m 0.1
a
f v
m 0.1
a
d 1 2 3 4


