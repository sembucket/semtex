#
# Example of a "script" for setting up an sview scene
#

f w
m 0.1
a
m -.1
t 0 0 0
p -135 155 0
z 1
d
